----------------------------------------------------------------------------------
-- Domipheus Labs - ArtyS7_RPU_SoC
--
-- SoC implementation for Digilent Arty S7-50. RPU rv32i RISV-V CPU, 192KB block ram
-- 256MB DDR3, SPI interface for SD card, and 720p HDMI/DVI-D textual output.
--
--
-- Tested with Vivado 2018.1
--
-- Author: Colin Riley
-- Twitter: @domipheus
--
-- Copyright 2018 Colin Riley
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

use IEEE.NUMERIC_STD.ALL;

library UNISIM;
use UNISIM.VComponents.all;

use work.constants.all;

entity rpu_top is
    Port ( 
    -- Input 100MHz clock
    CLK100MHZ : in STD_LOGIC;
    
    -- Input switches from board
    sw : in STD_LOGIC_VECTOR (3 downto 0);
    
    -- Output leds to board
    led : out STD_LOGIC_VECTOR (3 downto 0);
    	 
    -- SPI master interface 1
    O_spim1_sclk: out STD_LOGIC;
    I_spim1_miso: in STD_LOGIC;
    O_spim1_mosi: out STD_LOGIC;
    O_spim1_cs:   out STD_LOGIC;
    O_spim1_cd:   out STD_LOGIC;
    
    -- DDR3 interface
    ddr3_dq       : inout std_logic_vector(15 downto 0);
    ddr3_dqs_p    : inout std_logic_vector(1 downto 0);
    ddr3_dqs_n    : inout std_logic_vector(1 downto 0);

    ddr3_addr     : out   std_logic_vector(13 downto 0);
    ddr3_ba       : out   std_logic_vector(2 downto 0);
    ddr3_ras_n    : out   std_logic;
    ddr3_cas_n    : out   std_logic;
    ddr3_we_n     : out   std_logic;
    ddr3_reset_n  : out   std_logic;
    ddr3_ck_p     : out   std_logic_vector(0 downto 0);
    ddr3_ck_n     : out   std_logic_vector(0 downto 0);
    ddr3_cke      : out   std_logic_vector(0 downto 0);
    ddr3_cs_n     : out   std_logic_vector(0 downto 0);
    ddr3_dm       : out   std_logic_vector(1 downto 0);
    ddr3_odt      : out   std_logic_vector(0 downto 0);
    
    -- HDMI (DVI-D) video output
    hdmi_out_p : out STD_LOGIC_VECTOR(3 downto 0);
    hdmi_out_n : out STD_LOGIC_VECTOR(3 downto 0)
);
end rpu_top;

architecture Behavioral of rpu_top is
 
    -- DDR3 memory controller. This is generated by Xilinx MIG for 7-series FPGAs
    component mig_7series_0
        port(
            ddr3_dq       : inout std_logic_vector(15 downto 0);
            ddr3_dqs_p    : inout std_logic_vector(1 downto 0);
            ddr3_dqs_n    : inout std_logic_vector(1 downto 0);
            
            ddr3_addr     : out   std_logic_vector(13 downto 0);
            ddr3_ba       : out   std_logic_vector(2 downto 0);
            ddr3_ras_n    : out   std_logic;
            ddr3_cas_n    : out   std_logic;
            ddr3_we_n     : out   std_logic;
            ddr3_reset_n  : out   std_logic;
            ddr3_ck_p     : out   std_logic_vector(0 downto 0);
            ddr3_ck_n     : out   std_logic_vector(0 downto 0);
            ddr3_cke      : out   std_logic_vector(0 downto 0);
            ddr3_cs_n     : out   std_logic_vector(0 downto 0);
            ddr3_dm       : out   std_logic_vector(1 downto 0);
            ddr3_odt      : out   std_logic_vector(0 downto 0);
            
            app_addr                  : in    std_logic_vector(27 downto 0);
            app_cmd                   : in    std_logic_vector(2 downto 0);
            app_en                    : in    std_logic;
            app_wdf_data              : in    std_logic_vector(127 downto 0);
            app_wdf_end               : in    std_logic;
            app_wdf_mask              : in    std_logic_vector(15 downto 0);
            app_wdf_wren              : in    std_logic;
            app_rd_data               : out   std_logic_vector(127 downto 0);
            app_rd_data_end           : out   std_logic;
            app_rd_data_valid         : out   std_logic;
            app_rdy                   : out   std_logic;
            app_wdf_rdy               : out   std_logic;
            app_sr_req                : in    std_logic;
            app_ref_req               : in    std_logic;
            app_zq_req                : in    std_logic;
            app_sr_active             : out   std_logic;
            app_ref_ack               : out   std_logic;
            app_zq_ack                : out   std_logic;
            
            ui_clk                    : out   std_logic;
            ui_clk_sync_rst           : out   std_logic;
            init_calib_complete       : out   std_logic;
            -- System Clock Ports
            sys_clk_i                 : in    std_logic;
            -- Reference Clock Ports
            clk_ref_i       : in    std_logic;
            device_temp_i   : in    std_logic_vector(11 downto 0);
            device_temp     : out std_logic_vector(11 downto 0);
            sys_rst         : in std_logic
        );
    end component mig_7series_0;


    -- The RPU core definition
    COMPONENT core
        PORT(
            I_clk : IN  std_logic;
            I_reset : IN  std_logic;
            I_halt : IN  std_logic;
            I_int : IN  std_logic;
            O_int_ack : OUT  std_logic;
            
            MEM_O_cmd : OUT  std_logic;
            MEM_O_we : OUT  std_logic;
            
            MEM_O_byteEnable : OUT  std_logic_vector(1 downto 0);
            MEM_O_addr : OUT  std_logic_vector(31 downto 0);
            MEM_O_data : OUT  std_logic_vector(31 downto 0);
            MEM_I_data : IN  std_logic_vector(31 downto 0);
            
            MEM_I_ready : IN  std_logic;
            MEM_I_dataReady : IN  std_logic
            
            ;
            O_DBG:out std_logic_vector(XLEN32M1 downto 0)
        );
    END COMPONENT;
    
    COMPONENT clocking
        generic (
            in_mul    : natural := 10;    
            pix_div   : natural := 30;
            pix5x_div : natural := 10
        );
        PORT ( 
            I_unbuff_clk         : in  STD_LOGIC;
            O_buff_clkpixel      : out  STD_LOGIC;
            O_buff_clk5xpixel    : out  STD_LOGIC;
            O_buff_clk5xpixelinv : out  STD_LOGIC
        );
    END COMPONENT;
    
    
    -- This is generated by the Xilinx block ram generator
    -- Internally it simply utilizes multiple block ram primitives to give a view of a
    -- 64KB true dual-port ram device.
    component BRAM_64KB_wrapper is
        port (
            I_addra : in STD_LOGIC_VECTOR ( 31 downto 0 );
            I_clka : in STD_LOGIC;
            I_dina : in STD_LOGIC_VECTOR ( 31 downto 0 );
            O_douta : out STD_LOGIC_VECTOR ( 31 downto 0 );
            I_ena : in STD_LOGIC;
            I_wea : in STD_LOGIC_VECTOR ( 3 downto 0 );
            I_addrb : in STD_LOGIC_VECTOR ( 31 downto 0 );
            I_clkb : in STD_LOGIC;
            I_dinb : in STD_LOGIC_VECTOR ( 31 downto 0 );
            O_doutb : out STD_LOGIC_VECTOR ( 31 downto 0 );
            I_enb : in STD_LOGIC;
            I_web : in STD_LOGIC_VECTOR ( 3 downto 0 )
        );
    end component BRAM_64KB_wrapper;
    
    COMPONENT vga_gen
        generic (
            hRez       : natural := 1280;    
            hStartSync : natural := 1280+72;
            hEndSync   : natural := 1280+72+80;
            hMaxCount  : natural := 1280+72+80+216;
            hsyncActive : std_logic := '0';
            
            vRez       : natural := 720;
            vStartSync : natural := 720+3;
            vEndSync   : natural := 720+3+5;
            vMaxCount  : natural := 720+3+5+22;
            vsyncActive : std_logic := '1';
            prefetch_idx:natural := 8
        );
        PORT(    
            pixel_clock  : in std_logic; 
            pixel_h      : out STD_LOGIC_VECTOR(11 downto 0);
            pixel_v      : out STD_LOGIC_VECTOR(11 downto 0);
            pixel_h_pref : out STD_LOGIC_VECTOR(11 downto 0) := (others => '0');
            pixel_v_pref : out STD_LOGIC_VECTOR(11 downto 0) := (others => '0');
            blank_pref   : OUT std_logic;
            blank        : OUT std_logic;
            hsync        : OUT std_logic;
            vsync        : OUT std_logic
        );
    END COMPONENT;
    
    COMPONENT dvid
        PORT(
            clk      : IN std_logic;
            clk_n    : IN std_logic;
            clk_pixel: IN std_logic;
            red_p    : IN std_logic_vector(7 downto 0);
            green_p  : IN std_logic_vector(7 downto 0);
            blue_p   : IN std_logic_vector(7 downto 0);
            blank    : IN std_logic;
            hsync    : IN std_logic;
            vsync    : IN std_logic;          
            red_s    : OUT std_logic;
            green_s  : OUT std_logic;
            blue_s   : OUT std_logic;
            clock_s  : OUT std_logic
        );
    END COMPONENT;
    
    --- character generator
    
    
    COMPONENT char_generator is
        Port ( 
            I_clk_pixel : in  STD_LOGIC;
            
            -- Inputs from VGA signal generator
            -- defines the 'next pixel' 
            I_blank : in  STD_LOGIC;
            I_x : in  STD_LOGIC_VECTOR (11 downto 0);
            I_y : in  STD_LOGIC_VECTOR (11 downto 0);
            
            -- Request data for a glyph row from FRAM
            O_FRAM_ADDR : out STD_LOGIC_VECTOR (15 downto 0);
            I_FRAM_DATA : in STD_LOGIC_VECTOR (15 downto 0);
            
            -- Request data from textual memory TRAM
            O_TRAM_ADDR : out STD_LOGIC_VECTOR (15 downto 0);
            I_TRAM_DATA : in STD_LOGIC_VECTOR (15 downto 0);
            
            -- The data for the relevant requested pixel
            O_R : out STD_LOGIC_VECTOR (7 downto 0);
            O_G : out STD_LOGIC_VECTOR (7 downto 0);
            O_B : out STD_LOGIC_VECTOR (7 downto 0)
        );
    end COMPONENT;
    
    
    COMPONENT font_rom is
        port(
            clk: in std_logic;
            addr: in std_logic_vector(11 downto 0);
            data: out std_logic_vector(7 downto 0)
        );
    end COMPONENT;
     
    COMPONENT spi_master
        PORT(
            clock : IN  std_logic;
            reset_n : IN  std_logic;
            enable : IN  std_logic;
            cpol : IN  std_logic;
            cpha : IN  std_logic;
            cont : IN  std_logic;
            clk_div : IN integer;
            addr : IN  integer;
            tx_data : IN  std_logic_vector(7 downto 0);
            miso : IN  std_logic;
            sclk : buffer  std_logic;
            ss_n : buffer  std_logic_vector(7 downto 0);
            mosi : OUT  std_logic;
            busy : OUT  std_logic;
            rx_data : OUT  std_logic_vector(7 downto 0)
        );
    END COMPONENT;
        
    
    signal count: unsigned(31 downto 0) := X"00000000";
    
    -- Clock engine    
    signal cEng_pixel_720 : std_logic;
    signal cEng_5xpixel_720 : std_logic;    
    signal cEng_5xpixel_inv_720 : std_logic;
    
    -- Vga timing
    signal pixel_h : STD_LOGIC_VECTOR(11 downto 0);
    signal pixel_v : STD_LOGIC_VECTOR(11 downto 0);
    signal blank   : std_logic;
    signal hsync   : std_logic;
    signal vsync   : std_logic;    
    
    -- prefetch timing
    signal pixel_h_pref : STD_LOGIC_VECTOR(11 downto 0);
    signal pixel_v_pref : STD_LOGIC_VECTOR(11 downto 0);
    signal blank_pref: std_logic;
    
    signal	O_DBG: std_logic_vector(XLEN32M1 downto 0);
    
    signal cEng_core : std_logic := '0';
    signal I_reset : std_logic := '1';
    signal I_halt : std_logic := '0';
    signal I_int : std_logic := '0';
    signal MEM_I_ready : std_logic := '1';
    signal MEM_I_data : std_logic_vector(31 downto 0) := (others => '0');
    signal MEM_I_dataReady : std_logic := '0';



    signal MEM_O_data_swizzed : std_logic_vector(31 downto 0) := (others => '0');
 
 
    signal O_int_ack : std_logic;
    
    signal MEM_O_cmd : std_logic := '0';
    signal MEM_O_we : std_logic := '0';
    signal MEM_O_byteEnable : std_logic_vector(1 downto 0) := (others => '0');
    signal MEM_O_addr : std_logic_vector(31 downto 0) := (others => '0');
    signal MEM_O_data : std_logic_vector(31 downto 0) := (others => '0');


    signal mI_wea : STD_LOGIC_VECTOR ( 3 downto 0 ):= (others => '0');
    signal mI_clkb : STD_LOGIC;
    signal mI_dinb : STD_LOGIC_VECTOR ( 31 downto 0 ):= (others => '0');
    signal mO_doutb : STD_LOGIC_VECTOR ( 31 downto 0 ):= (others => '0');
    signal mI_enb : STD_LOGIC;
    signal mI_web : STD_LOGIC_VECTOR ( 3 downto 0 );
    signal mI_enb_others_0 : STD_LOGIC:= '0';

    -- Clock period definitions
    constant I_clk_period : time := 3 ns;
    
    
    signal IO_LEDS: STD_LOGIC_VECTOR(7 downto 0):= (others => '0');
    signal INT_DATA: std_logic_vector(BWIDTHM1 downto 0):= (others => '0');
    signal IO_DATA: std_logic_vector(BWIDTHM1 downto 0):= (others => '0');
    signal DDR3_DATA: std_logic_vector(BWIDTHM1 downto 0):= (others => '0');
    
    -- Block ram management
    signal MEM_64KB_ADDR : std_logic_vector(31 downto 0):= (others => '0');
    signal MEM_BANK_ID : std_logic_vector(15 downto 0):= (others => '0');
    signal MEM_ANY_CS : std_logic := '0';
    signal MEM_WE : std_logic := '0';
    
    signal MEM_CS_BRAM_1 : std_logic := '0';
    signal MEM_CS_BRAM_2 : std_logic := '0';
    signal MEM_CS_BRAM_3 : std_logic := '0';
    
    
    signal MEM_CS_DDR3 : std_logic := '0';
    
    signal MEM_CS_SYSTEM : std_logic := '0';
    
    signal MEM_DATA_OUT_BRAM_1: std_logic_vector(BWIDTHM1 downto 0):= (others => '0');
    signal MEM_DATA_OUT_BRAM_2: std_logic_vector(BWIDTHM1 downto 0):= (others => '0');
    signal MEM_DATA_OUT_BRAM_3: std_logic_vector(BWIDTHM1 downto 0):= (others => '0');
   
    signal red_s   : std_logic:= '0';
    signal green_s : std_logic:= '0';
    signal blue_s  : std_logic:= '0';
    signal clock_s : std_logic:= '0';
    
    ----------------------------------------------------------------------------
    -- Text Graphics Subsystem
    
    signal SYS_TRAM1_OUTDATA: std_logic_vector(15 downto 0);
    signal SYS_TRAM2_OUTDATA: std_logic_vector(15 downto 0);
    signal SYS_TRAM_2K_ADDR: std_logic_vector(15 downto 0);
    
    signal SYS_FRAM1_ADDR: std_logic_vector(15 downto 0);
    signal SYS_FRAM1_OUTDATA: std_logic_vector(15 downto 0);
    
    signal SYS_FRAM2_ADDR: std_logic_vector(15 downto 0);
    signal SYS_FRAM2_OUTDATA: std_logic_vector(15 downto 0);
    
    
    signal GFX_MODE: std_logic := '0';  -- 0 = text 1 = pixel
    
    signal TXT_R: std_logic_vector(7 downto 0);
    signal TXT_G: std_logic_vector(7 downto 0);
    signal TXT_B: std_logic_vector(7 downto 0);
    
    signal FRAM_DATA: std_logic_vector(15 downto 0);
    signal FRAM_ADDR: std_logic_vector(15 downto 0);
    
    
    signal FRAM_DATA_TEST: std_logic_vector(7 downto 0);
    signal FRAM_ADDR_TEST: std_logic_vector(11 downto 0);
    
    signal TRAM_DATA: std_logic_vector(15 downto 0);
    signal TRAM_ADDR: std_logic_vector(15 downto 0);
    
    signal tram_32b_addr : STD_LOGIC_VECTOR ( 31 downto 0 ):= (others => '0');
    
    
    signal MEM_I_data_raw : std_logic_vector(31 downto 0) := (others => '0');
    
    
    --Inputs
    signal spim1_clock : std_logic := '0';
    signal spim1_reset_n : std_logic := '1';
    signal spim1_enable : std_logic := '0';
    signal spim1_cpol : std_logic := '0';
    signal spim1_cpha : std_logic := '0';
    signal spim1_cont : std_logic := '0';
    signal spim1_clk_div : integer := 10;
    signal spim1_addr : integer:= 0;
    signal spim1_tx_data : std_logic_vector(7 downto 0) := (others => '0');
    signal spim1_miso : std_logic := '1';
    
    --Outputs
    signal spim1_sclk : std_logic:='0';
    signal spim1_ss_n : std_logic_vector(1 downto 0):= (others => '1');
    signal spim1_mosi : std_logic;
    signal spim1_busy : std_logic := '0';
    signal spim1_rx_data : std_logic_vector(7 downto 0);

    constant ADDR_WIDTH            : integer := 28;

    signal init_calib_complete_i       : std_logic:= '0';
    signal device_temp                 : std_logic_vector(11 downto 0):= (others => '1'); 
    signal app_addr                    : std_logic_vector(27 downto 0):= (others => '1');
    signal app_addr_i                  : std_logic_vector(31 downto 0):= (others => '1');
    signal app_cmd                     : std_logic_vector(2 downto 0):= (others => '1');
    signal app_en                      : std_logic:= '0';
    signal app_rdy                     : std_logic:= '0';
    signal app_rdy_i                   : std_logic:= '0';
    signal app_rd_data                 : std_logic_vector(127 downto 0):= (others => '1');
    signal app_rd_data_end             : std_logic:= '0';
    signal app_rd_data_valid           : std_logic:= '0';
    signal app_rd_data_valid_i         : std_logic:= '0';
    signal app_wdf_data                : std_logic_vector(127 downto 0):= (others => '1');
    signal app_wdf_end                 : std_logic:= '1';
    signal app_wdf_mask                : std_logic_vector(15 downto 0):= (others => '0');
    signal app_wdf_rdy                 : std_logic:= '0';
    signal app_wdf_rdy_i               : std_logic:= '0';
    signal app_sr_active               : std_logic:= '0';
    signal app_ref_ack                 : std_logic:= '0';
    signal app_zq_ack                  : std_logic:= '0';
    signal app_wdf_wren                : std_logic:= '0';
    
    signal device_temp_i                 :    std_logic_vector(11 downto 0):= (others => '1');
    signal clk                         : std_logic:= '0';
    signal rst                         : std_logic:= '0';
    signal sys_rst                     :     std_logic:= '0';
    
    signal ddr3_sys_clk_i :     std_logic:= '0';
    signal ddr3_clk_ref_i :     std_logic:= '0';
    
    
    signal ddr3_rd_buffer                : std_logic_vector(127 downto 0):= (others => '0');
    
    
    -- UI app clock output from MIG
    signal ddr3_ui_clk: std_logic:= '0';
    signal ddr3_ui_clk_unbuff: std_logic:= '0';
    signal Clk_Mem: std_logic:= '0';
    signal Clk_Soc: std_logic:= '0';
    
    
    constant MIG_DDR3_CMD_WRITE: std_logic_vector(2 downto 0) := "000";
    constant MIG_DDR3_CMD_READ: std_logic_vector(2 downto 0) := "001";
    
    signal memcontroller_ddr3_state: integer := 0;
    
    -- Documentation says to giv
    signal memcontroller_reset_count: integer := 100000;
    
    signal CLK200MHZ: std_logic := '0';
    

    type ddr3_mask_lookup_t is array (0 to 3) of std_logic_vector(3 downto 0);
    
    constant ddr3_16b_wmask : ddr3_mask_lookup_t := 
    ( "0011",
      "0011",
      "1100",
      "1100" );
    
    constant ddr3_8b_wmask : ddr3_mask_lookup_t := 
    ( "0111",
      "1011",
      "1101",
      "1110" );

    --- PERFORMANCE COUNTERS
    signal counter_clock_cycles_core : std_logic_vector(31 downto 0) := X"00000000";
    signal counter_clock_cycles_core_last_calc : std_logic_vector(31 downto 0) := X"00000000";
    signal counter_clock_cycles_mem : std_logic_vector(31 downto 0) := X"00000000";
    signal counter_clock_cycles_mem_last_calc : std_logic_vector(31 downto 0) := X"00000000";
    signal counter_clock_cycles_soc : std_logic_vector(31 downto 0) := X"00000000";
    signal counter_clock_cycles_soc_last_calc : std_logic_vector(31 downto 0) := X"00000000";
    
    signal counter_clock_cycles_100mhz : std_logic_vector(31 downto 0) := X"00000000";
    signal counter_clock_cycles_100mhz_secondcount : std_logic_vector(31 downto 0) := X"00000000"; 
    
    signal counter_clock_freq_core : std_logic_vector(31 downto 0) :=   X"00000000";
    signal counter_clock_freq_mem : std_logic_vector(31 downto 0) := X"00000000";
    signal counter_clock_freq_soc : std_logic_vector(31 downto 0) := X"00000000";
    
    signal counter_ddr3_read_req  : std_logic_vector(31 downto 0) := X"00000000";
    signal counter_ddr3_write_req  : std_logic_vector(31 downto 0) := X"00000000";
    signal counter_ddr3_cmdready_read_wait_cycles  : std_logic_vector(31 downto 0) := X"00000000";
    signal counter_ddr3_read_wait_cycles  : std_logic_vector(31 downto 0) := X"00000000";
    signal counter_ddr3_cmdready_write_wait_cycles  : std_logic_vector(31 downto 0) := X"00000000";
    signal counter_ddr3_write_wait_cycles  : std_logic_vector(31 downto 0) := X"00000000";


    signal MEM_readyState: integer := 0;
    signal MEM_readyState_stable:integer := 0;
    signal DDR3_ReadyState: integer := 0;
    signal DDR3_ReadyState_stable:integer := 0;
    
    -- DDR3_CtrState definitions - running off MEM clock domain
    constant DDR3_CtlState_Ready : integer :=  0;
    constant DDR3_CtlState_ReadCmdIssued : integer :=   1;
    constant DDR3_CtlState_ReadCmdComplete: integer  :=   2;
    constant DDR3_CtlState_WriteCmdIssued : integer  :=  5;
    constant DDR3_CtlState_WriteCmdComplete : integer  :=  6;
    
    -- SOC_CtrState definitions - running off SOC clock domain
    constant SOC_CtlState_Ready : integer :=  0;
    
    -- IMM SOC control states are immediate 1-cycle latency
    -- i.e. BRAM or explicit IO
    constant SOC_CtlState_IMM_WriteCmdComplete : integer := 9;
    constant SOC_CtlState_IMM_ReadCmdComplete : integer := 6;
    
    -- DDR3 SOC control states have unknown latency and cross clock domains.
    -- SOC_* and DDR3*_ state flags are used as flags to sync valid data
    -- across the different clocked domains.
    constant SOC_CtlState_DDR3_ReadCmdIssued : integer := 10;
    constant SOC_CtlState_DDR3_ReadCmdInFlight : integer := 11;
    constant SOC_CtlState_DDR3_ReadCmdComplete: integer  := 12;
    constant SOC_CtlState_DDR3_WriteCmdIssued : integer  := 20;
    constant SOC_CtlState_DDR3_WriteCmdInFlight : integer  := 21;
    constant SOC_CtlState_DDR3_WriteCmdComplete : integer  := 22;


    function F_ChangeEndian ( data : in std_logic_vector ) return std_logic_vector  is
        constant numBytes: integer := data'length/8;
    begin
        assert(numBytes = 4);
        return data(7 downto 0) & data(15 downto 8) & data(23 downto 16) & data(31 downto 24);
    end function F_ChangeEndian; 

BEGIN

    ddr3_init_waiter: process(CLK100MHZ)
    begin
        if rising_edge(CLK100MHZ) then
            if (memcontroller_reset_count > 0) then
                memcontroller_reset_count <= memcontroller_reset_count - 1;
            end if;
        end if;
    end process;
    
    -- The DDR3 reset is held active low at the start, and the CPU
    -- reset is held active high for the same amount of time.
    sys_rst <= '1' when (memcontroller_reset_count = 0) else '0';
    I_reset <= '0' when (memcontroller_reset_count = 0) else '1';

    clk_core_count: process(cEng_core)
    begin
        if rising_edge(cEng_core) then
            counter_clock_cycles_core <= std_logic_vector(unsigned(counter_clock_cycles_core) + 1);
        end if;
    end process;
        
    Clk_Mem_count: process(Clk_Mem)
    begin
        if rising_edge(Clk_Mem) then
           counter_clock_cycles_mem <= std_logic_vector(unsigned(counter_clock_cycles_mem) + 1);
        end if;
    end process;
    
    Clk_Soc_count: process(cEng_core)
    begin
        if rising_edge(cEng_core) then
          counter_clock_cycles_soc <= std_logic_vector(unsigned(counter_clock_cycles_soc) + 1);
        end if;
    end process;
    
    -- increment the counter each 100MHz cycle
    process(CLK100MHZ)
    begin
        if rising_edge(CLK100MHZ) then
            count <= count + 1;
        end if;
    end process;
        
    clk_100mhz_count: process(CLK100MHZ)
    begin
       if rising_edge(CLK100MHZ) then
           counter_clock_cycles_100mhz <= std_logic_vector(unsigned(counter_clock_cycles_100mhz) + 1);
           
           if counter_clock_cycles_100mhz_secondcount = X"05f5e100" then -- 100,000,000
              counter_clock_cycles_100mhz_secondcount <= X"00000000";
              counter_clock_freq_core <= std_logic_vector(unsigned(counter_clock_cycles_core) - unsigned(counter_clock_cycles_core_last_calc));
              counter_clock_freq_soc <= std_logic_vector(unsigned(counter_clock_cycles_soc) - unsigned(counter_clock_cycles_soc_last_calc));
              counter_clock_freq_mem <= std_logic_vector(unsigned(counter_clock_cycles_mem) - unsigned(counter_clock_cycles_mem_last_calc));
           else
              counter_clock_cycles_100mhz_secondcount <= std_logic_vector(unsigned(counter_clock_cycles_100mhz_secondcount) + 1);
              
              if counter_clock_cycles_100mhz_secondcount = X"00000001" then
                counter_clock_cycles_core_last_calc <= counter_clock_cycles_core;
                counter_clock_cycles_mem_last_calc <= counter_clock_cycles_mem;
                counter_clock_cycles_soc_last_calc <= counter_clock_cycles_soc;
              end if;
           end if;   
       end if;
    end process;

    -- Move MEM_readyState into the Clk_Mem domain *_stable
    MEM_readyState_TryStable : process(Clk_Mem)
    begin
        if rising_edge(Clk_Mem) then
            MEM_readyState_stable <= MEM_readyState;
        end if;
    end process;
    
    -- Move DDR3_ReadyState into the Clk_Soc/Core domain *_stable
    DDR3_ReadyState_TryStable : process(cEng_core)
    begin
        if rising_edge(cEng_core) then
            DDR3_ReadyState_stable <= DDR3_ReadyState;
        end if;
    end process;

 -- DDR3 memory interface. Generated using Xilinx Memory Interface Generator.
 u_mig_7series_0 : mig_7series_0
      port map (
       -- Memory interface ports
       ddr3_addr                      => ddr3_addr,
       ddr3_ba                        => ddr3_ba,
       ddr3_cas_n                     => ddr3_cas_n,
       ddr3_ck_n                      => ddr3_ck_n,
       ddr3_ck_p                      => ddr3_ck_p,
       ddr3_cke                       => ddr3_cke,
       ddr3_ras_n                     => ddr3_ras_n,
       ddr3_reset_n                   => ddr3_reset_n,
       ddr3_we_n                      => ddr3_we_n,
       ddr3_dq                        => ddr3_dq,
       ddr3_dqs_n                     => ddr3_dqs_n,
       ddr3_dqs_p                     => ddr3_dqs_p,
       init_calib_complete            => init_calib_complete_i,
       device_temp                    => device_temp,
       ddr3_cs_n                      => ddr3_cs_n,
       ddr3_dm                        => ddr3_dm,
       ddr3_odt                       => ddr3_odt,
-- Application interface ports
       app_addr                       => app_addr,
       app_cmd                        => app_cmd,
       app_en                         => app_en,
       app_wdf_data                   => app_wdf_data,
       app_wdf_end                    => app_wdf_end,
       app_wdf_wren                   => app_wdf_wren,
       app_rd_data                    => app_rd_data,
       app_rd_data_end                => app_rd_data_end,
       app_rd_data_valid              => app_rd_data_valid,
       app_rdy                        => app_rdy,
       app_wdf_rdy                    => app_wdf_rdy,
       app_sr_req                     => '0',
       app_ref_req                    => '0',
       app_zq_req                     => '0',
       app_sr_active                  => app_sr_active,
       app_ref_ack                    => app_ref_ack,
       app_zq_ack                     => app_zq_ack,
       ui_clk                         => Clk_Mem, --ddr3_ui_clk,
       ui_clk_sync_rst                => rst,
       app_wdf_mask                   => app_wdf_mask,
-- System Clock Ports
       sys_clk_i                      => CLK100MHZ,
-- Reference Clock Ports
       clk_ref_i                      => CLK200MHZ,
       device_temp_i                  => device_temp_i,
       sys_rst                        => sys_rst
        );
-- End of User Design top instance
 
 	-- The O_we signal can sustain too long. Clamp it to only when O_cmd is active.
    MEM_WE <= MEM_O_cmd and MEM_O_we;
    
    -- "Local" BRAM banks are 64KB. To address inside we need lower 16b
    MEM_64KB_ADDR <= X"0000" & MEM_O_addr(15 downto 0);
    MEM_BANK_ID <= MEM_O_addr(31 downto 16);

    MEM_CS_BRAM_1 <= '1' when (MEM_BANK_ID = X"0000") else '0'; -- 0x0000ffff bank 64KB
    MEM_CS_BRAM_2 <= '1' when (MEM_BANK_ID = X"0001") else '0'; -- 0x0001ffff bank 64KB
    MEM_CS_BRAM_3 <= '1' when (MEM_BANK_ID = X"0002") else '0'; -- 0x0002ffff bank 64KB
    
    MEM_CS_DDR3 <= '1' when (MEM_BANK_ID(15 downto 12) = X"1") else '0'; -- 0x1******* ddr3 bank 256MB
    
    -- if any CS line is active, this is 1
    MEM_ANY_CS <= MEM_CS_BRAM_1 or MEM_CS_BRAM_2 or MEM_CS_BRAM_3;
    
    -- select the correct data to send to cpu
    MEM_I_data_raw <= INT_DATA when O_int_ack = '1'     
                  else MEM_DATA_OUT_BRAM_1 when MEM_CS_BRAM_1 = '1' 
                  else MEM_DATA_OUT_BRAM_2 when MEM_CS_BRAM_2 = '1' 
                  else MEM_DATA_OUT_BRAM_3 when MEM_CS_BRAM_3 = '1' 
                  else IO_DATA;
 
    -- Endian swizzles occuring here on the falling edges of clocks.
    -- This should be moved into the CPU core.
    data_in_endian_swizz: process(cEng_core)
    begin 
        if falling_edge(cEng_core) then
            case MEM_O_byteEnable is
               when "10" =>
                
                    MEM_I_data <=   MEM_I_data_raw( 7 downto 0) & MEM_I_data_raw(15 downto 8) & MEM_I_data_raw(23 downto 16) & MEM_I_data_raw(31 downto 24);
               when "01" =>
                  
                        case MEM_O_addr(1 downto 0) is
                            when "00" =>
                              -- unaligned...
                              MEM_I_data <= X"0000" & MEM_I_data_raw(23 downto 16) & MEM_I_data_raw(31 downto 24);
                            when "01" =>
                              MEM_I_data <= X"0000" & MEM_I_data_raw(23 downto 16) & MEM_I_data_raw(31 downto 24);
                            when "10" =>
                              -- unaligned...
                              MEM_I_data <= X"0000" & MEM_I_data_raw( 7 downto 0) & MEM_I_data_raw(15 downto 8);
                            when "11" =>
                              MEM_I_data <= X"0000" & MEM_I_data_raw( 7 downto 0) & MEM_I_data_raw(15 downto 8);
                            when others =>
                        end case;
                    
               when "00" =>

                    case MEM_O_addr(1 downto 0) is
                        when "00" =>
                            MEM_I_data <= X"000000" & MEM_I_data_raw(31 downto 24);
                        when "01" =>
                            MEM_I_data <= X"000000" & MEM_I_data_raw(23 downto 16);
                        when "10" =>
                            MEM_I_data <= X"000000" & MEM_I_data_raw(15 downto 8);
                        when "11" =>
                            MEM_I_data <= X"000000" & MEM_I_data_raw( 7 downto 0);
                        when others =>
                    end case;
                when others =>
            end case;
        end if;
    end process;
    
    data_out_endian_swizz: process(cEng_core)
    begin 
        if falling_edge(cEng_core) then
        if (MEM_WE = '1') then
            case MEM_O_byteEnable is
               when "10" =>
                    mI_wea <= "1111";
                  
                  MEM_O_data_swizzed <= MEM_O_data( 7 downto 0) & MEM_O_data(15 downto 8) & MEM_O_data(23 downto 16) & MEM_O_data(31 downto 24);
               when "01" =>
                    case MEM_O_addr(1 downto 0) is
                        
                        when "00" =>
                          mI_wea <= "1100";
                          MEM_O_data_swizzed <=  MEM_O_data( 7 downto 0) & MEM_O_data(15 downto 8) & X"0000" ;
                        when "01" =>
                           --  unaligned
                          mI_wea <= "1100";
                          MEM_O_data_swizzed <= MEM_O_data( 7 downto 0) & MEM_O_data(15 downto 8) & X"0000" ;
                        when "10" =>
                          mI_wea <= "0011";
                          MEM_O_data_swizzed <= X"0000" & MEM_O_data( 7 downto 0) & MEM_O_data(15 downto 8);
                        when "11" =>
                          --this is unaligned, shouldn't be supported...
                          mI_wea <= "0011";
                          MEM_O_data_swizzed <=  X"0000" & MEM_O_data( 7 downto 0) & MEM_O_data(15 downto 8);
                        when others =>
                    end case;
               when "00" =>

                     case MEM_O_addr(1 downto 0) is
                           when "00" =>
                               mI_wea <= "1000";
                             MEM_O_data_swizzed <=  MEM_O_data(7 downto 0) & X"000000";
                           when "01" =>
                               mI_wea <= "0100";
                             MEM_O_data_swizzed <= X"00" & MEM_O_data(7 downto 0) & X"0000"; 
                           when "10" =>
                               mI_wea <= "0010";
                             MEM_O_data_swizzed <=  X"0000" & MEM_O_data( 7 downto 0) & X"00";
                           when "11" =>
                               mI_wea <= "0001";
                             MEM_O_data_swizzed <= X"000000" & MEM_O_data( 7 downto 0);
                           when others =>
                       end case;
                when others =>
            end case;
            else

            mI_wea <= "0000";
            end if;
        end if;
    end process;
    
    
    spi_m_1: spi_master PORT MAP (            
         clock => cEng_core, 
         reset_n => spim1_reset_n,            
         enable => spim1_enable, 
         cpol => spim1_cpol,
         cpha => spim1_cpha,
         cont => spim1_cont,
         clk_div => spim1_clk_div,
         addr => spim1_addr,
         tx_data => spim1_tx_data,
         miso => spim1_miso,
         sclk => spim1_sclk,
         mosi => spim1_mosi,
         busy => spim1_busy,
         rx_data => spim1_rx_data
       );
       
       O_spim1_cd <= '0';
       O_spim1_sclk <=spim1_sclk;
       spim1_miso <= I_spim1_miso;
       O_spim1_mosi <= spim1_mosi;
       O_spim1_cs <= spim1_ss_n(1);
       
       clkEngine_200: clocking
       generic map (
           in_mul  => 10,
           pix_div => 5,
           pix5x_div => 7
       )
       port map (
           I_unbuff_clk => CLK100MHZ,
           O_buff_clkpixel => CLK200MHZ, 
           O_buff_clk5xpixel => cEng_core,
           O_buff_clk5xpixelinv => open
       ); 


   core0: core PORT MAP (
          I_clk => cEng_core,
          I_reset => I_reset,
          I_halt => I_halt,
          I_int => I_int,
          O_int_ack => O_int_ack,
          MEM_I_ready => MEM_I_ready,
          MEM_O_cmd => MEM_O_cmd,
          MEM_O_we => MEM_O_we,
          MEM_O_byteEnable => MEM_O_byteEnable,
          MEM_O_addr => MEM_O_addr,
          MEM_O_data => MEM_O_data,
          MEM_I_data => MEM_I_data,
          MEM_I_dataReady => MEM_I_dataReady
		  ,
		  O_DBG=>O_DBG
        );
        
   mem1: BRAM_64KB_wrapper port map (
       I_addra => MEM_64KB_ADDR,
       I_clka => cEng_core,
       I_dina => MEM_O_data_swizzed,
       O_douta => MEM_DATA_OUT_BRAM_1,
       I_ena => MEM_CS_BRAM_1,
       I_wea => mI_wea,
       I_addrb => tram_32b_addr,
       I_clkb => cEng_pixel_720,
       I_dinb => mI_dinb,
       O_doutb => open,
       I_enb => mI_enb,
       I_web => mI_web
   );     
   
   mem2: BRAM_64KB_wrapper port map (
       I_addra => MEM_64KB_ADDR,
       I_clka => cEng_core,
       I_dina => MEM_O_data_swizzed,
       O_douta => MEM_DATA_OUT_BRAM_2,
       I_ena => MEM_CS_BRAM_2,
       I_wea => mI_wea,
       I_addrb => tram_32b_addr,
       I_clkb => cEng_pixel_720,
       I_dinb => mI_dinb,
       O_doutb => mO_doutb,
       I_enb => mI_enb,
       I_web => mI_web
   ); 
          
   mem3: BRAM_64KB_wrapper port map (
      I_addra => MEM_64KB_ADDR,
      I_clka => cEng_core,
      I_dina => MEM_O_data_swizzed,
      O_douta => MEM_DATA_OUT_BRAM_3,
      I_ena => MEM_CS_BRAM_3,
      I_wea => mI_wea,
      I_addrb => tram_32b_addr,
      I_clkb => cEng_pixel_720,
      I_dinb => mI_dinb,
      O_doutb => open,
      I_enb => mI_enb,
      I_web => mI_web
      );


    -- Huge process which handles memory request arbitration at the Soc/Core clock 
    MEM_proc: process(cEng_core)
    begin
        if rising_edge(cEng_core) then
            if MEM_readyState = SOC_CtlState_Ready then
                if MEM_O_cmd = '1' then
                
                    -- system memory maps
                    if MEM_O_addr = X"f0009000" and MEM_O_we = '1' then
                        -- onboard leds
                        IO_LEDS <= "0000" & MEM_O_data( 3 downto 0);
                    end if;

                    -- spi -- needs adjusted for endian
                    if MEM_O_addr = X"f0009300" and MEM_O_we = '1' then
                        spim1_reset_n <= MEM_O_data_swizzed(27); --LSB[3]
                        spim1_cpol <= MEM_O_data_swizzed(26); --LSB[2]
                        spim1_cpha <= MEM_O_data_swizzed(25); --LSB[1]
                        spim1_cont <= MEM_O_data_swizzed(24); --LSB[0]
                    end if;
                    
                    if MEM_O_addr = X"f000930c" and MEM_O_we = '1' then
                        spim1_clk_div <= to_integer(unsigned( std_logic_vector'( (MEM_O_data_swizzed(23 downto 16)) & (MEM_O_data_swizzed(31 downto 24))))) ;
                    end if;
                    
                    if MEM_O_addr = X"f000930e" and MEM_O_we = '1' then
                        spim1_addr <= to_integer(unsigned(MEM_O_data_swizzed(26 downto 24)));
                        -- raw CS line select
                        spim1_ss_n(1) <= MEM_O_data_swizzed(24); 
                    end if;
                    
                    -- spi -- needs adjusted for endian
                    if MEM_O_addr = X"f0009300" and MEM_O_we = '0' then
                        IO_DATA(31 downto 28) <= "0000";
                        IO_DATA(27) <= spim1_reset_n;
                        IO_DATA(26) <= spim1_cpol;
                        IO_DATA(25) <= spim1_cpha;
                        IO_DATA(24) <= spim1_cont;
                        IO_DATA(23 downto 8) <= std_logic_vector(to_unsigned(spim1_clk_div, 16));
                        IO_DATA(7 downto 3) <= "00000";
                        IO_DATA(2 downto 0) <= "00" & spim1_ss_n(1);--std_logic_vector(to_unsigned(spim1_addr, 3));
            
                    end if;
                    
                    if MEM_O_addr = X"f0009304" and MEM_O_we = '0' then
                       --little endian
                       IO_DATA(31 downto 0) <= X"0" & "000" & spim1_busy & X"000000" ;
                    
                    end if;
                     
                    if MEM_O_addr = X"f0009308" and MEM_O_we = '0' then
                       --little endian
                       IO_DATA(31 downto 0) <= spim1_rx_data & X"000000";
                    end if;
                    
                    if MEM_O_addr = X"f0009308" and MEM_O_we = '1' and spim1_busy = '0' then
                        spim1_tx_data <= MEM_O_data_swizzed(31 downto 24); -- LSByte
                        spim1_enable <= '1';
                    end if;
                    
                    -- DDR3 config registers
                    if MEM_O_addr = X"fdd30000" and MEM_O_we = '0' then
                        --little endian
                        IO_DATA(31 downto 0) <= "0000000" & init_calib_complete_i & X"000000";
                    end if;
                    
                    -- perf counters
                    
                   if MEM_O_addr = X"ff001000" and MEM_O_we = '0' then
                     IO_DATA <= F_ChangeEndian(counter_clock_cycles_core);
                   end if; 
                        
                   if MEM_O_addr = X"ff001004" and MEM_O_we = '0' then
                     IO_DATA <= F_ChangeEndian(counter_clock_cycles_100mhz);
                   end if;
                   
                   if MEM_O_addr = X"ff001008" and MEM_O_we = '0' then
                     IO_DATA <= F_ChangeEndian(counter_clock_freq_core);
                   end if;
                   
                   if MEM_O_addr = X"ff00100C" and MEM_O_we = '0' then
                     IO_DATA <= F_ChangeEndian(counter_clock_freq_mem);
                   end if;
                                        
                    if MEM_O_addr = X"ff001010" and MEM_O_we = '0' then
                      IO_DATA <= F_ChangeEndian(counter_clock_freq_soc);
                    end if;
                  
                   if MEM_O_addr = X"ff001100" and MEM_O_we = '0' then
                     IO_DATA <= F_ChangeEndian(counter_ddr3_read_req);
                   end if;
                   
                   if MEM_O_addr = X"ff001104" and MEM_O_we = '0' then
                     IO_DATA <= F_ChangeEndian(counter_ddr3_write_req);
                   end if;
                   
                   if MEM_O_addr = X"ff001108" and MEM_O_we = '0' then
                     IO_DATA <= F_ChangeEndian(counter_ddr3_cmdready_read_wait_cycles);
                   end if;
                   
                   if MEM_O_addr = X"ff00110c" and MEM_O_we = '0' then
                     IO_DATA <= F_ChangeEndian(counter_ddr3_read_wait_cycles);
                   end if;
                    
                    if MEM_O_addr = X"ff001110" and MEM_O_we = '0' then
                      IO_DATA <= F_ChangeEndian(counter_ddr3_cmdready_write_wait_cycles);
                    end if;
                   
                   if MEM_O_addr = X"ff001114" and MEM_O_we = '0' then
                     IO_DATA <= F_ChangeEndian(counter_ddr3_write_wait_cycles);
                   end if;
                   
                   
                    -- DDR3 burst read debug reading
                    if MEM_O_addr = X"ffff0000" and MEM_O_we = '0' then
                         IO_DATA <= ddr3_rd_buffer(127 downto 96);
                    end if;
                    if MEM_O_addr = X"ffff0004" and MEM_O_we = '0' then
                        IO_DATA <= ddr3_rd_buffer(95 downto 64);
                    end if;
                    if MEM_O_addr = X"ffff0008" and MEM_O_we = '0' then
                       IO_DATA <= ddr3_rd_buffer(63 downto 32);
                    end if;
                    if MEM_O_addr = X"ffff000c" and MEM_O_we = '0' then
                       IO_DATA <= ddr3_rd_buffer(31 downto 0);
                    end if;
                    
                    -- DDR3 burst write debug reading
                    if MEM_O_addr = X"ffff0010" and MEM_O_we = '0' then
                         IO_DATA <= app_wdf_data(127 downto 96);
                    end if;
                    if MEM_O_addr = X"ffff0014" and MEM_O_we = '0' then
                        IO_DATA <= app_wdf_data(95 downto 64);
                    end if;
                    if MEM_O_addr = X"ffff0018" and MEM_O_we = '0' then
                       IO_DATA <= app_wdf_data(63 downto 32);
                    end if;
                    if MEM_O_addr = X"ffff001c" and MEM_O_we = '0' then
                       IO_DATA <= app_wdf_data(31 downto 0);
                    end if;
                    
                    MEM_I_ready <= '0';
                    MEM_I_dataReady  <= '0';
                    if MEM_O_we = '1' then
                        -- DDR3 request, or immediate command?
                        if MEM_CS_DDR3 = '1' then
                           MEM_readyState <= SOC_CtlState_DDR3_WriteCmdIssued;
                           counter_ddr3_write_req <= std_logic_vector(unsigned(counter_ddr3_write_req) + 1);
                        else
                           MEM_readyState <= SOC_CtlState_IMM_WriteCmdComplete;
                        end if;
                    else
                        -- DDR3 request, or immediate command?
                        if MEM_CS_DDR3 = '1' then
                            MEM_readyState <= SOC_CtlState_DDR3_ReadCmdIssued;
                            counter_ddr3_read_req <= std_logic_vector(unsigned(counter_ddr3_read_req) + 1);
                        else
                            MEM_readyState <= SOC_CtlState_IMM_ReadCmdComplete;
                        end if;
                    end if;
                    
                end if;
            elsif MEM_readyState >= 1 then
                
                spim1_enable <= '0';
                
                -- Immediate commands do not cross clock domains and complete immediately
                if MEM_readyState = SOC_CtlState_IMM_ReadCmdComplete then
                    MEM_I_ready <= '1';
                    MEM_I_dataReady <= '1'; 
                    MEM_readyState <= SOC_CtlState_Ready;  
                    
                elsif MEM_readyState = SOC_CtlState_IMM_WriteCmdComplete then
                    MEM_I_ready <= '1';
                    MEM_I_dataReady  <= '0'; 
                    MEM_readyState <= SOC_CtlState_Ready;
                    
                -- DDR3 read states ****(crosses clock domain)****
                elsif MEM_readyState = SOC_CtlState_DDR3_ReadCmdIssued then
                    if (DDR3_ReadyState_stable = DDR3_CtlState_ReadCmdIssued) then
                        MEM_readyState <= SOC_CtlState_DDR3_ReadCmdInFlight;
                    end if;
                elsif MEM_readyState = SOC_CtlState_DDR3_ReadCmdInFlight then    
                    if DDR3_ReadyState_stable = DDR3_CtlState_ReadCmdComplete then
                        MEM_readyState <= SOC_CtlState_DDR3_ReadCmdComplete;
                    end if;
                elsif MEM_readyState = SOC_CtlState_DDR3_ReadCmdComplete then    
                    IO_DATA <= DDR3_DATA;
                    MEM_I_ready <= '1';
                    MEM_I_dataReady <= '1'; 
                    MEM_readyState <= SOC_CtlState_Ready; 
                    
                   
                -- DDR3 write states ****(crosses clock domain)****            
                elsif MEM_readyState = SOC_CtlState_DDR3_WriteCmdIssued then
                    if DDR3_ReadyState_stable = DDR3_CtlState_WriteCmdIssued then
                        MEM_readyState <= SOC_CtlState_DDR3_WriteCmdInFlight;
                    end if;
                elsif MEM_readyState = SOC_CtlState_DDR3_WriteCmdInFlight then   
                    if DDR3_ReadyState_stable = DDR3_CtlState_WriteCmdComplete then
                        MEM_readyState <= SOC_CtlState_DDR3_WriteCmdComplete;
                    end if;
                elsif MEM_readyState = SOC_CtlState_DDR3_WriteCmdComplete then
                    MEM_I_ready <= '1';
                    MEM_I_dataReady  <= '0'; 
                    MEM_readyState <= SOC_CtlState_Ready;
                    
                else
                    MEM_readyState <= MEM_readyState + 1;
                end if;
            end if;
        end if;
    end process;

    -- DDR3 Request handler, runs at Memory clock.
    -- Needs to read data across the SOC clock domain.
    DDR3_proc: process(Clk_Mem)
    begin
        if rising_edge(Clk_Mem) then
            if DDR3_ReadyState = DDR3_CtlState_Ready then
                if MEM_readyState_stable = SOC_CtlState_DDR3_WriteCmdIssued  then
                    -- DDR3 Write
                    if app_rdy = '1' and app_wdf_rdy = '1' then                 
                          app_addr <= '0' & MEM_O_addr(27 downto 1);
                          app_cmd <= MIG_DDR3_CMD_WRITE;
                          app_en <= '1';
                          
                          app_wdf_wren <= '1';
                          
                          case MEM_O_byteEnable is
                              when "10" =>
                                  if MEM_O_addr(3 downto 2) = "00" then
                                      app_wdf_data <= MEM_O_data_swizzed & X"AAAAAAAA" & X"BBBBBBBB" & X"CCCCCCCC";
                                      app_wdf_mask <= X"0FFF";
                                  elsif MEM_O_addr(3 downto 2) = "01" then
                                      app_wdf_data <= X"AAAAAAAA" & MEM_O_data_swizzed & X"BBBBBBBB" & X"CCCCCCCC";
                                      app_wdf_mask <= X"F0FF";
                                  elsif MEM_O_addr(3 downto 2) = "10" then
                                      app_wdf_data <= X"AAAAAAAA" & X"BBBBBBBB" & MEM_O_data_swizzed & X"CCCCCCCC";
                                      app_wdf_mask <= X"FF0F";
                                  elsif MEM_O_addr(3 downto 2) = "11" then
                                      app_wdf_data <= X"AAAAAAAA" & X"BBBBBBBB" & X"CCCCCCCC" & MEM_O_data_swizzed;
                                      app_wdf_mask <= X"FFF0";
                                  end if; 
                              when "01" =>
                                  if MEM_O_addr(3 downto 2) = "00" then
                                      app_wdf_data <= MEM_O_data_swizzed & X"AAAAAAAA" & X"BBBBBBBB" & X"CCCCCCCC";
                                      app_wdf_mask <= ddr3_16b_wmask(to_integer(unsigned(MEM_O_addr(1 downto 0)))) & X"FFF";
                                  elsif MEM_O_addr(3 downto 2) = "01" then
                                      app_wdf_data <= X"AAAAAAAA" & MEM_O_data_swizzed & X"BBBBBBBB" & X"CCCCCCCC";
                                      app_wdf_mask <= X"F" & ddr3_16b_wmask(to_integer(unsigned(MEM_O_addr(1 downto 0)))) & X"FF";
                                  elsif MEM_O_addr(3 downto 2) = "10" then
                                      app_wdf_data <= X"AAAAAAAA" & X"BBBBBBBB" & MEM_O_data_swizzed & X"CCCCCCCC";
                                      app_wdf_mask <= X"FF" & ddr3_16b_wmask(to_integer(unsigned(MEM_O_addr(1 downto 0)))) & X"F";
                                  elsif MEM_O_addr(3 downto 2) = "11" then
                                      app_wdf_data <= X"AAAAAAAA" & X"BBBBBBBB" & X"CCCCCCCC" & MEM_O_data_swizzed;
                                      app_wdf_mask <= X"FFF" & ddr3_16b_wmask(to_integer(unsigned(MEM_O_addr(1 downto 0))));
                                  end if; 
                             when "00" =>
                                 if MEM_O_addr(3 downto 2) = "00" then
                                     app_wdf_data <= MEM_O_data_swizzed & X"AAAAAAAA" & X"BBBBBBBB" & X"CCCCCCCC";
                                     app_wdf_mask <= ddr3_8b_wmask(to_integer(unsigned(MEM_O_addr(1 downto 0)))) & X"FFF";
                                 elsif MEM_O_addr(3 downto 2) = "01" then
                                     app_wdf_data <= X"AAAAAAAA" & MEM_O_data_swizzed & X"BBBBBBBB" & X"CCCCCCCC";
                                     app_wdf_mask <= X"F" & ddr3_8b_wmask(to_integer(unsigned(MEM_O_addr(1 downto 0)))) & X"FF";
                                 elsif MEM_O_addr(3 downto 2) = "10" then
                                     app_wdf_data <= X"AAAAAAAA" & X"BBBBBBBB" & MEM_O_data_swizzed & X"CCCCCCCC";
                                     app_wdf_mask <= X"FF" & ddr3_8b_wmask(to_integer(unsigned(MEM_O_addr(1 downto 0)))) & X"F";
                                 elsif MEM_O_addr(3 downto 2) = "11" then
                                     app_wdf_data <= X"AAAAAAAA" & X"BBBBBBBB" & X"CCCCCCCC" & MEM_O_data_swizzed;
                                     app_wdf_mask <= X"FFF" & ddr3_8b_wmask(to_integer(unsigned(MEM_O_addr(1 downto 0))));
                                 end if;
                              when others =>
                          end case;
                          DDR3_ReadyState <= DDR3_CtlState_WriteCmdIssued;
                        else
                          counter_ddr3_cmdready_write_wait_cycles <= std_logic_vector(unsigned(counter_ddr3_cmdready_write_wait_cycles) + 1);                
                      end if;  
                      
                elsif MEM_readyState_stable = SOC_CtlState_DDR3_ReadCmdIssued  then
                    -- DDR3 Read
                    if app_rdy = '1' then
                      app_addr <= '0' &  MEM_O_addr(27 downto 1);
                      app_cmd <= MIG_DDR3_CMD_READ;
                      app_en <= '1';
                      DDR3_ReadyState <= DDR3_CtlState_ReadCmdIssued;
                    else
                       counter_ddr3_cmdready_read_wait_cycles <= std_logic_vector(unsigned(counter_ddr3_cmdready_read_wait_cycles) + 1);
                    end if;
                end if;
            elsif DDR3_ReadyState = DDR3_CtlState_ReadCmdIssued then
                   if app_rdy = '1' and app_en = '1' then
                     app_en <= '0';
                   end if;
          
                   if app_rd_data_valid = '1' then
                      ddr3_rd_buffer <= app_rd_data;
                      case MEM_O_byteEnable is
                          when "10" =>
                               DDR3_DATA(31 downto 0) <= app_rd_data(127 downto 96);
                          when "01" =>
                               case MEM_O_addr(1 downto 0) is
                                  when "00" =>
                                    DDR3_DATA(31 downto 0) <= app_rd_data(127 downto 112) & X"AAAA";
                                  when "01" =>
                                    DDR3_DATA(31 downto 0) <= app_rd_data(127 downto 112) & X"BBBB";
                                  when "10" =>
                                    DDR3_DATA(31 downto 0) <= X"AAAA" & app_rd_data(95 downto 80);
                                  when "11" =>
                                     DDR3_DATA(31 downto 0) <= X"BBBB" & app_rd_data(95 downto 80);
                                  when others =>
                              end case;
                               
                          when "00" =>                              
                                case MEM_O_addr(1 downto 0) is
                               when "00" => 
                                      DDR3_DATA(31 downto 0) <= app_rd_data(127 downto 120) & X"AAAAAA"; 
                                    when "01" =>
                                      DDR3_DATA(31 downto 0) <=  X"BB" &app_rd_data(119 downto 112) & X"BBBB"; 
                                    when "10" =>
                                      DDR3_DATA(31 downto 0) <= X"CCCC" & app_rd_data(95 downto 88) & X"CC"; 
                                    when "11" =>
                                      DDR3_DATA(31 downto 0) <= X"DDDDDD" & app_rd_data(87 downto 80); 
                                    when others =>
                                end case;
                          when others =>
                      end case;

                      DDR3_ReadyState <= DDR3_CtlState_ReadCmdComplete;
                  else
                     counter_ddr3_read_wait_cycles <= std_logic_vector(unsigned(counter_ddr3_read_wait_cycles) + 1); 
                  end if;
            elsif DDR3_ReadyState = DDR3_CtlState_ReadCmdComplete then
              if MEM_readyState_stable = SOC_CtlState_Ready then
                DDR3_ReadyState <= DDR3_CtlState_Ready;
              end if;  
            elsif DDR3_ReadyState = DDR3_CtlState_WriteCmdIssued then
                 if app_rdy = '1' and app_en = '1' then
                   app_en <= '0';
                 end if;
         
                 if app_wdf_rdy = '1' and app_wdf_wren = '1' then
                   app_wdf_wren <= '0';
                 end if;
                 
                if MEM_readyState_stable = SOC_CtlState_DDR3_WriteCmdInFlight  then
                     if app_en = '0' and app_wdf_wren = '0' then
                         DDR3_ReadyState <= DDR3_CtlState_WriteCmdComplete;
                     end if;
                end if;
                 counter_ddr3_write_wait_cycles <= std_logic_vector(unsigned(counter_ddr3_write_wait_cycles) + 1);   
                 
            elsif DDR3_ReadyState = DDR3_CtlState_WriteCmdComplete then
                 if MEM_readyState_stable = SOC_CtlState_Ready then
                   DDR3_ReadyState <= DDR3_CtlState_Ready;
                 end if;  
            end if;
        end if;
    end process;


   -- Gen 75Mhz pixel clock generation
   -- Technically, 720p should be 74.25MHz. 75 generally works on monitors. YMMV.
   clock_eng_1280_720A: clocking
    generic map (
        in_mul  => 9,
        pix_div => 12,
        pix5x_div => 12
    )
    port map (
        I_unbuff_clk => CLK100MHZ,
        O_buff_clkpixel => cEng_pixel_720,
        O_buff_clk5xpixel => open,
        O_buff_clk5xpixelinv => open
    );   
    
   clock_eng_1280_720B: clocking
   generic map (
       in_mul  => 10,
       pix_div => 1,
       pix5x_div => 2
   )
   port map (
       I_unbuff_clk => cEng_pixel_720,
       O_buff_clkpixel => open,
       O_buff_clk5xpixel => cEng_5xpixel_720,
       O_buff_clk5xpixelinv => cEng_5xpixel_inv_720
   );   
    
    Inst_vga_gen: vga_gen 
    generic map (
        hRez        => 1280,
        hStartSync  => 1280+72,
        hEndSync    => 1280+72+80,
        hMaxCount   => 1280+72+80+216,
        hsyncActive => '0',
        vRez        => 720,
        vStartSync  => 720+3,
        vEndSync    => 720+3+5,
        vMaxCount   => 720+3+5+22,
        vsyncActive => '1'
    )
    PORT MAP( 
        pixel_clock  => cEng_pixel_720,    
        pixel_h      => pixel_h,
        pixel_v      => pixel_v,
        pixel_h_pref => pixel_h_pref,
        pixel_v_pref => pixel_v_pref,     
        blank_pref   => blank_pref,
        blank        => blank,
        hsync        => hsync,
        vsync        => vsync
    );
            
    -- at the moment I'm using an external font rom and the above frams
    -- are not connected This will change in the future, so glyphs can be dynamically
    -- altered with different fonts
    fram_test: 
    font_rom port map(
       clk => cEng_pixel_720,
       addr => FRAM_ADDR_TEST,
       data => FRAM_DATA_TEST
    );
    
    FRAM_ADDR_TEST <= FRAM_ADDR(11 downto 0);
    FRAM_DATA <= X"00" & FRAM_DATA_TEST;
       
    text_generator_engine: char_generator PORT MAP (
        I_clk_pixel => cEng_pixel_720,
        
        I_blank => blank_pref,
        I_x => pixel_h_pref ,
        I_y => pixel_v_pref ,
        
        O_FRAM_ADDR => FRAM_ADDR,
        I_FRAM_DATA => FRAM_DATA,
        
        O_TRAM_ADDR => TRAM_ADDR,
        I_TRAM_DATA => TRAM_DATA,
        
        O_R => TXT_R,
        O_G => TXT_G, 
        O_B => TXT_B
    );
       
    -- Tram uses 16 bit addressing
    -- just address the 32 bit of our block ram, data will be swizzled automatically.
    tram_32b_addr <= X"0000" & TRAM_ADDR(15 downto 0);   
    mI_enb <= '1';
    mI_web <= "0000";
            
    -- Select the 16 bits required
    TRAM_DATA <= mO_doutb(31 downto 24)& mO_doutb(23 downto 16)  when (TRAM_ADDR(1) = '0') else  mO_doutb(15 downto 8) &  mO_doutb(7 downto 0);
    
    -- TMDS signal generation
    -- This takes pixel colour values and synd data, generating the
    -- 10-bit coding.
    dvid_1: dvid PORT MAP(
        clk        => cEng_5xpixel_720,
        clk_n      => cEng_5xpixel_inv_720, 
        clk_pixel  => cEng_pixel_720,
        red_p      => TXT_R,
        green_p    => TXT_G,
        blue_p     => TXT_B,
        blank      => blank,
        hsync      => hsync,
        vsync      => vsync,
        
        -- outputs to TMDS drivers
        red_s      => red_s,
        green_s    => green_s,
        blue_s     => blue_s,
        clock_s    => clock_s
    );
    
	OBUFDS_blue  : OBUFDS port map ( O  => hdmi_out_p(0), OB => hdmi_out_n(0), I  => blue_s );
	OBUFDS_green   : OBUFDS port map ( O  => hdmi_out_p(1), OB => hdmi_out_n(1), I  => green_s );
	OBUFDS_red : OBUFDS port map ( O  => hdmi_out_p(2), OB => hdmi_out_n(2), I  => red_s );
	OBUFDS_clock : OBUFDS port map ( O  => hdmi_out_p(3), OB => hdmi_out_n(3), I  => clock_s );

    led <= IO_LEDS(3 downto 0); 
end Behavioral;
